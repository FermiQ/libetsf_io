netcdf read_dim_t01 {
dimensions:
	number_of_atom_species = 2 ;
	number_of_atoms = 5 ;
	character_string_length = 80 ;
	number_of_reduced_dimensions = 3 ;
	number_of_vectors = 3 ;
variables:
	char atom_species_names(number_of_atom_species, character_string_length) ;
	int atom_species(number_of_atoms) ;
	double reduced_atom_positions(number_of_atoms, number_of_reduced_dimensions) ;
	double primitive_vectors(number_of_vectors, number_of_reduced_dimensions) ;

// global attributes:
		:file_format = "ETSF Nanoquanta" ;
		:file_format_version = 1.3f ;
		:Conventions = "http://www.etsf.eu/fileformats" ;
		:title = "Silane molecule generated by ncgen." ;
data:

 atom_species_names =
  "Si",
  "H" ;

 atom_species = 1, 2, 2, 2, 2 ;

 reduced_atom_positions =
  0.5, 0.5, 0.5,
  0.6, 0.6, 0.6,
  0.4, 0.4, 0.6,
  0.6, 0.4, 0.4,
  0.4, 0.6, 0.4 ;

 primitive_vectors =
  10, 0, 0,
  0, 10, 0,
  0, 0, 10 ;
}
