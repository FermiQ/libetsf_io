netcdf test_write_electrons {
dimensions:
	character_string_length = 80 ;
	max_number_of_angular_momenta = 1 ;
	max_number_of_coefficients = 6 ;
	max_number_of_projectors = 2 ;
	max_number_of_states = 8 ;
	number_of_atoms = 4 ;
	number_of_atom_species = 1 ;
	number_of_cartesian_directions = 3 ;
	number_of_components = 2 ;
	number_of_grid_points_vector1 = 1 ;
	number_of_grid_points_vector2 = 1 ;
	number_of_grid_points_vector3 = 5 ;
	number_of_kpoints = 12 ;
	my_number_of_kpoints = 6;
	number_of_reduced_dimensions = 3 ;
	number_of_spinor_components = 1 ;
	number_of_spins = 1 ;
	number_of_symmetry_operations = 4 ;
	number_of_vectors = 3 ;
	real_or_complex = 1 ;
	symbol_length = 2 ;
variables:
	int my_kpoints(my_number_of_kpoints);
	int number_of_electrons ;
	char exchange_functional(character_string_length) ;
	char correlation_functional(character_string_length) ;
	double fermi_energy ;
		fermi_energy:units = "Klingon units" ;
		fermi_energy:scale_to_atomic_units = 0.123 ;
	char smearing_scheme(character_string_length) ;
	double smearing_width ;
		smearing_width:units = "atomic units" ;
		smearing_width:scale_to_atomic_units = 1. ;
	int number_of_states(number_of_spins, my_number_of_kpoints) ;
	double eigenvalues(number_of_spins, my_number_of_kpoints, max_number_of_states) ;
		eigenvalues:units = "atomic units" ;
		eigenvalues:scale_to_atomic_units = 1. ;
	double occupations(number_of_spins, my_number_of_kpoints, max_number_of_states) ;

// global attributes:
		:file_format = "ETSF Nanoquanta" ;
		:file_format_version = 1.3f ;
		:Conventions = "http://www.etsf.eu/fileformats/" ;
		:title = "Test" ;
		:history = "" ;
data:

 number_of_electrons = 1 ;

 exchange_functional = "aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa" ;

 correlation_functional = "aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa" ;

 fermi_energy = 1 ;

 smearing_scheme = "aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa" ;

 smearing_width = 1 ;

 my_kpoints =
  1, 3, 5, 7, 11, 12 ;

 number_of_states =
  1, 3, 5, 7, 11, 12 ;

 eigenvalues =
  1, 2, 3, 4, 5, 6, 7, 8,
  17, 18, 19, 20, 21, 22, 23, 24,
  33, 34, 35, 36, 37, 38, 39, 40,
  49, 50, 51, 52, 53, 54, 55, 56,
  81, 82, 83, 84, 85, 86, 87, 88,
  89, 90, 91, 92, 93, 94, 95, 96 ;

 occupations =
  1, 2, 3, 4, 5, 6, 7, 8,
  17, 18, 19, 20, 21, 22, 23, 24,
  33, 34, 35, 36, 37, 38, 39, 40,
  49, 50, 51, 52, 53, 54, 55, 56,
  81, 82, 83, 84, 85, 86, 87, 88,
  89, 90, 91, 92, 93, 94, 95, 96 ;
}
