netcdf Test {
dimensions:
  number_of_atom_species = 2;
  number_of_atoms = 5;
  character_string_length = 80;
  number_of_reduced_dimensions = 3;
  number_of_vectors = 3;
  number_of_components = 2;

variables:
  char atom_species_names(number_of_atom_species, character_string_length);
  int atom_species(number_of_atoms);
  int test_integer_2d(number_of_atom_species, number_of_atom_species);
  int test_integer_4d(number_of_components, number_of_vectors, number_of_vectors, number_of_atom_species);
  int space_group;
  double test_double_0d;
  double test_double_1d(number_of_vectors);
  double reduced_atom_positions(number_of_atoms, number_of_reduced_dimensions);
  double primitive_vectors(number_of_vectors, number_of_reduced_dimensions);
  double density(number_of_components, number_of_vectors, number_of_vectors, number_of_vectors);

  // Global attributes
  :file_format = "ETSF Nanoquanta";
  :file_format_version = 1.3f;
  :Conventions = "http://www.etsf.eu/fileformats";
  :title = "Silane molecule generated by ncgen.";

data:
  space_group = 1;
  atom_species_names = "Si", "H";
  atom_species = 1, 2, 2, 2, 2;
  test_integer_2d = 1, 2, 3, 4;
  test_integer_4d = 1, 2, 3, 4, 5, 6, 7, 8, 9,
                    10, 11, 12, 13, 14, 15, 16, 17, 18,
                    -1, -2, -3, -4, -5, -6, -7, -8, -9,
                    -10, -11, -12, -13, -14, -15, -16, -17, -18;
  test_double_0d = 3.14;
  test_double_1d = 1., 2., 3.;
  reduced_atom_positions = 0.5, 0.5, 0.5, 0.6, 0.6, 0.6, 0.4, 0.4, 0.6, 0.6, 0.4, 0.4, 0.4, 0.6, 0.4;
  primitive_vectors = 10., 0., 0., 0., 10., 0., 0., 0., 10.;
  density = 0., 1., 0., 1., 2., 1., 0., 1., 0.,
            1., 2., 1., 2., 3., 2., 1., 2., 1.,
            0., 1., 0., 1., 2., 1., 0., 1., 0.,
            -0., -1., -0., -1., -2., -1., -0., -1., -0.,
            -1., -2., -1., -2., -3., -2., -1., -2., -1.,
            -0., -1., -0., -1., -2., -1., -0., -1., -0.;
}
